module inst_mem(  
    input clk, reset, 
    input [31:0] pc,  
    output reg [31:0] instruction  
    );  
    wire [3:0] rom_addr = pc[9:2];  
    reg [31:0] rom[255:0];  // 256 words of 32 bits each
    initial begin  
//---------------------------------------------Different Type Instruction-----------------------------------------------------------------        
//        rom[0] = 32'b001000_00000_00001_0000000000000100; // addi $s1, $s0, 4
//        rom[1] = 32'b001000_00001_00010_0000000000000010; // addi $s2, $s1, 2
//        rom[2] = 32'b000000_00000_00001_00011_00000_100000; // add $s3, $s0, $s1
//        rom[3] = 32'b000000_00010_00001_00011_00000_100100; // and $s3, $s2, $s1
//        rom[4] = 32'b101011_00010_00011_0000000000001000; // sw $s3, $s2, 8
//        rom[5] = 32'b100011_00010_00100_0000000000010000; // lw $s4, $s2, 16
//        rom[6] = 32'b100011_10011_00101_0000000000010000; // lw $s5, $s2, 16
//        rom[7] = 32'b00010010001100100000000000010000; // beq $s1, $s2, 4
//        rom[8] = 32'b00100010000101010000000000000100; // addi $s1, $s0, 4
//        rom[9] = 32'b00001000000000000000000000000101; // j 5
//        rom[10] = 32'b00000000000000000000000000000000; // nop
//        rom[11] = 32'b00000000000000000000000000000000; // nop
//        rom[12] = 32'b00000000000000000000000000000000; // nop
//---------------------------------------------One Clock Cycle Hazard -----------------------------------------------------------------       
//        rom[0] = 32'b001000_00000_00001_0000000000000001; // addi $1, $0, 1
//        rom[1] = 32'b001000_00001_00011_0000000000000011; // addi $3, $1, 3
//        rom[2] = 32'b001000_00000_00101_0000000000000101; // addi $5 $0, 5
//        // EX_MEM Rd  ID_EX Rs Hazard  --> $2
//        rom[3] = 32'b00000_00001_00011_00010_00000_100000; //add $2,   $1, $3
//        rom[4] = 32'b00000_00010_00101_01100_00000_100100; //and $12, $2, $5
//        rom[5] = 32'b00000000000000000000000000000000; // nop
//        rom[6] = 32'b00000000000000000000000000000000; // nop
//        rom[7] = 32'b00000000000000000000000000000000; // nop        
        // EX_MEM Rd  ID_EX Rt Hazard  --> $2
//        rom[0] = 32'b00000_00001_00011_00010_00000_100000; //add $2,   $1, $3
//        rom[1] = 32'b00000_00101_00010_01100_00000_100100; //and $12, $5, $2
//---------------------------------------------Two Clock Cycle Hazard -----------------------------------------------------------------           
////        // MEM_WB Rd  ID_EX Rs Hazard  --> $2 <---Two Clock Cycle
//        rom[0] = 32'b00000_00001_00011_00010_00000_100000; //add $2,   $1, $3
//        rom[1] = 32'b00000_00101_00100_01100_00000_100100; //and $12, $5, $4
//        rom[2] = 32'b00000_00010_00110_01101_00000_100101; //or   $13, $2, $6
        
        // MEM_WB Rd   ID_EX Rs Hazard  --> $2 <---Two Clock Cycle
//        rom[0] = 32'b00000_00001_00011_00010_00000_100000; //add $2,   $1, $3
//        rom[1] = 32'b00000_00101_00010_00010_00000_100100; //and $2, $5, $2
//        rom[2] = 32'b00000_00110_00010_01101_00000_100101; //or   $13, $6 $2
//---------------------------------------------Test B-Type -----------------------------------------------------------------               
        rom[0] = 32'b000100_00000_00000_0000000000000010; // beq $s0, $0, 2
        rom[1] = 32'b00000_00101_00001_00011_00000_100100; //and $3, $5, $1
        rom[2] = 32'b00000_00110_00011_01101_00000_100101; //or   $13, $6 $3
        rom[3] = 32'b00000_00111_00011_01101_00000_100010; //sub   $13, $7 $3
        rom[4] = 32'b00000_01000_00011_01101_00000_100000; //add   $13, $8 $3
//---------------------------------------------Test Load Use Hazard-----------------------------------------------------------------           
//        rom[0] = 32'b100011_00001_00010_0000000000000000; // lw $2 , 0($1)  
//        rom[1] = 32'b000000_00010_00001_01100_00000_100100; // and $12, $2, $1
//        rom[2] = 32'b000000_00010_00001_01100_00000_100101; // or $12 $2 $1
//        rom[3] = 32'b00000000000000000000000000000000; // nop
//        rom[4] = 32'b00000000000000000000000000000000; // nop
    end  

    always@(*) begin
        if(reset)
            instruction =  32'd0;
        else
            instruction = (pc[31:0] < 32*8 )? rom[rom_addr]: 32'd0; 
    end
        
 endmodule   